`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:38:49 09/11/2018
// Design Name:   mux2
// Module Name:   U:/UB/Digital Logic and Design/Verilog/Lab2-1-New/Lab2-1-New/mux2_tb.v
// Project Name:  Lab2-1-New
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: mux2
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module mux2_tb;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	mux2 uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

